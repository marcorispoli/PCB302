********************************************************************************
* SN74HCS365.cir
* 2.0
* 2020-04-16 00:00:00
* Texas Instruments Incorporated.
* Standard Logic, SLHR
* 12500 TI Blvd
* Dallas, TX -75243
*
*
* Revision History:
* Rev 2.0: 01/01/2020
* - Model generated from datasheet values
* - Built using generic logic gate behavioral pspice model V2
* - Built using an automated model which generalizes parts under same family
* - Performance is expected typical behavior at 25C
* - Written for and tested with Tina-TI Version 9.3.100.244 SF-TI
* - Accurate power consumption with dyanmic as well as static Icc
*
********************************************************************************
*[Disclaimer]
* This model is designed as an aid for customers of Texas Instruments.
* TI and its licensors and suppliers make no warranties, either expressed
* or implied, with respect to this  model, including the warranties of
* merchantability or fitness for a particular purpose. The model is
* provided solely on an "as is" basis. The entire risk as to its quality
* and performance is with the customer.
*
*[Copyright]
*(C) Copyright 2020 Texas Instruments Incorporated. All rights reserved.
*
**
********************************************************************************
*                                 SN74HCS365
********************************************************************************
**1*.SUBCKT SN74HCS365 Y A VCC AGND

.SUBCKT SN74HCS365 Y A OEZ VCC AGND
XU1 Y A VCC OEZ VCC AGND LOGIC_GATE_2PIN_TRI_STATE_HC_1i_AND_Tristate_ST
.ENDS




*$
.SUBCKT LOGIC_GATE_2PIN_TRI_STATE_HC_1i_AND_Tristate_ST OUT A B OEZ VCC GND

.PARAM VCC_ABS_MAX = 7
.PARAM VCC_MAX = 6
.PARAM RA = 240000000
.PARAM RB = 240000000
.PARAM CA = 5e-12
.PARAM CB = 5e-12
.PARAM ROEZ = 5000
.PARAM COEZ = 3e-12
RA  A  GND {RA}
RB  B  GND {RB}
CA  A  GND {CA}
CB  B  GND {CB}
ROEZ OEZ GND {ROEZ}
COEZ OEZ GND {COEZ}
XUA NA A VCC GND LOGIC_INPUT_HC_1i_AND_Tristate_ST
XUB NB B VCC GND LOGIC_INPUT_HC_1i_AND_Tristate_ST
XUOEZ NOEZ OEZ VCC GND LOGIC_INPUT_HC_1i_AND_Tristate_ST
XUG NA NB NOUTG VCC GND LOGIC_FUNCTION_2_HC_1i_AND_Tristate_ST
XOUTPD NOUTG NOUTTPD VCC GND TPD_HC_1i_AND_Tristate_ST
XUOUT NOUTTPD NOUT_INT NOEZ VCC GND LOGIC_TRI_STATE_OUTPUT_HC_1i_AND_Tristate_ST
XICC VCC GND NVIOUT LOGIC_ICC_HC_1i_AND_Tristate_ST
SICC VCC GND VCC GND SW1
* Monitor Output Current *
H1 NVIOUT GND VIOUT 1 
VIOUT NOUT_INT OUTsw 0 
SIOFF OUTsw OUT VCC GND SW2
DA2 GND A D1
DB2 GND B D1
DO2 GND OUT D1
RDA1 NA1 GND 1e6 
RDB1 NB1 GND 1e6 
RDO1 NO1 GND 1e6 
DOE1 NOEZ VCC D1
DOE2 GND OEZ D1
SDA1 NA1 A VCC GND SW2
SDB1 NB1 B VCC GND SW2
SDO1 NO1 OUT VCC GND SW2
.MODEL SW1 VSWITCH VON = {VCC_ABS_MAX} VOFF = {VCC_MAX} RON = 10 ROFF = 60e6
.MODEL SW2 VSWITCH VON = {0.55} VOFF = {0.45} RON = 10m ROFF = 100e6
.MODEL D1 D
.ENDS
*$
.SUBCKT LOGIC_INPUT_HC_1i_AND_Tristate_ST OUT IN VCC VEE
.PARAM STANDARD_INPUT_SELECT = 0

.PARAM SCHMITT_TRIGGER_INPUT_SELECT = 1
ESTD_THR VSTD_THR VEE TABLE {V(VCC,VEE)} =
+(1,0.5)
+(1.8,0.9)
+(2.5,1.25)
+(3.3,1.65)
+(5,2.5)
+(6,3)
ETRP_P VTRP_P VEE TABLE {V(VCC,VEE)} =
+(2,1.2)
+(4.5,2.5)
+(6,3.3)
ETRP_N VTRP_N VEE TABLE {V(VCC,VEE)} =
+(2,0.6)
+(4.5,1.6)
+(6,2)
EHYST VHYST VEE TABLE {V(VCC,VEE)} =
+(2,0.6)
+(4.5,0.9)
+(6,1.3)
ETRUE NTRUE VEE VALUE = {V(VCC,VEE)}
EFALSE NFALSE VEE VALUE = {0}

EBETA BETA VEE VALUE = {V(VHYST,VEE)/(V(NTRUE,VEE) - V(NFALSE,VEE) + V(VHYST,VEE))}
EFB NFB VEE VALUE = {(1 - V(BETA,VEE))*V(IN,VEE) + V(BETA,VEE)*V(CURR_OUT,VEE)}
*EFB NFB VEE VALUE = {(1 - V(BETA,VEE))*V(IN,VEE) + V(BETA,VEE)*V(OUT,VEE)}
EREF NREF VEE VALUE = {0.5*(1 - V(BETA,VEE))*(V(VTRP_P,VEE) + V(VTRP_N,VEE)) 
+ + 0.5*V(BETA,VEE)*(V(NTRUE,VEE) + V(NFALSE,VEE))}
EDIFF NDIFF VEE VALUE = {V(NFB,NREF)}
*ECOMP OUT VEE VALUE = {0.5*V(VCC,VEE)*(SGN(V(NDIFF,VEE)) + ABS(SGN(V(NDIFF,VEE))))}
ESWITCH VSWITCH VEE VALUE = {0.5*(-SGN(V(NDIFF,VEE)) + ABS(SGN(V(NDIFF,VEE))))}
ESWITCH1 VSWITCH1 VEE VALUE = {0.5*(SGN(V(NDIFF,VEE)) + ABS(SGN(V(NDIFF,VEE))))}
GCOMP VEE CURR_OUT VALUE = {SCHMITT_TRIGGER_INPUT_SELECT*0.5*V(VCC,VEE)*(SGN(V(NDIFF,VEE)) + ABS(SGN(V(NDIFF,VEE))))}

GSTD VEE CURR_OUT VALUE = {STANDARD_INPUT_SELECT*0.5*V(VCC,VEE)*(SGN(V(IN,VSTD_THR)) + ABS(SGN(V(IN,VSTD_THR))))}
ROUT CURR_OUT VEE 1
EMID MID VEE VALUE = {0.5*(V(VCC,VEE) + V(VEE))}
EARG NARG VEE VALUE = {V(CURR_OUT,VEE) - V(MID,VEE)}
EOUT OUT VEE VALUE = {0.5*(SGN(V(NARG,VEE)) + ABS(SGN(V(NARG,VEE) ) ) )}
*EOUT OUT VEE CURR_OUT VEE 1

.PARAM MAXICC = .0009
.PARAM VT = .7
.PARAM VCC_MIN = 3

EV_VT1 VTN VEE VALUE = { VT }
EV_VT2 VTP VEE VALUE = { V(VCC,VEE) - VT }

ETEST TEST VEE VALUE = {.9*V(VCC,VEE)}

EVTHDIFF VTH_DIFF VEE VALUE = {V(IN,VSTD_THR)}
EVTHPDIFF VTHP_DIFF VEE VALUE = {V(IN,VTRP_P)}
EVTHNDIFF VTHN_DIFF VEE VALUE = {V(IN,VTRP_N)}
EVTNDIFF VTN_DIFF VEE VALUE = { V(IN,VTN) }
EVTPDIFF VTP_DIFF VEE VALUE = { V(IN,VTP) }


GICCVA VCC VEE VALUE = { (-ABS(( (1+SGN(V(VTN_DIFF,VEE)) ) )/2 -1) * 2*MAXICC*((V(IN,VEE)-VT)/V(VCC,VEE))^2)*(1 + SGN(V(VCC,VEE) - VCC_MIN))*V(VSWITCH,VEE)}
GICCVB VCC VEE VALUE = { (ABS(( (1+SGN(V(VTHP_DIFF,VEE)) ) )/2 -1) * 2*MAXICC*((V(IN,VEE)-VT)/V(VCC,VEE))^2)*(1 + SGN(V(VCC,VEE) - VCC_MIN))*V(VSWITCH,VEE)}

GICCVC VCC VEE VALUE = { ( ABS(  (1+SGN(V(VTHN_DIFF,VEE)) ) )/2     * 2*MAXICC*((V(IN,VEE)-(V(VCC,VEE)-VT))/V(VCC,VEE))^2)*(1 + SGN(V(VCC,VEE) - VCC_MIN))*V(VSWITCH1,VEE)}
GICCVD VCC VEE VALUE = { (-ABS(  (1+SGN(V(VTP_DIFF,VEE)) ) )/2     * 2*MAXICC*((V(IN,VEE)-(V(VCC,VEE)-VT))/V(VCC,VEE))^2)*(1 + SGN(V(VCC,VEE) - VCC_MIN))*V(VSWITCH1,VEE)}

.ENDS
*$
.SUBCKT LOGIC_FUNCTION_2_HC_1i_AND_Tristate_ST A B OUT VCC VEE
.PARAM AND  = 1
.PARAM NAND = 0
.PARAM OR   = 0
.PARAM NOR  = 0
.PARAM XOR  = 0
.PARAM XNOR = 0
GAND  VEE N1 VALUE = {AND*V(A,VEE)*V(B,VEE)}
GNAND VEE N1 VALUE = {NAND*(1 - V(A,VEE)*V(B,VEE))}
GOR   VEE N1 VALUE = {OR*(MIN(V(A,VEE) + V(B,VEE),1))}
GNOR  VEE N1 VALUE = {NOR*(1 - MIN(V(A,VEE) + V(B,VEE),1))}
GXOR  VEE N1 VALUE = {XOR*((1 - V(A,VEE))*V(B,VEE) + V(A,VEE)*(1 - V(B,VEE)))}
GXNOR VEE N1 VALUE = {XNOR*(1 - ((1 - V(A,VEE))*V(B,VEE) + V(A,VEE)*(1 - V(B,VEE))))}
RN1 N1 VEE 1
EOUT OUT VEE N1 VEE 1
.ENDS
*$
*$
.SUBCKT  TPD_HC_1i_AND_Tristate_ST IN OUT VCC VEE
.PARAM TPDELAY1 = 1N
.PARAM RS = 10K
.PARAM CS = {-TPDELAY1/(RS*LOG(0.5))}
*ETPDNORM NTPDNORM VEE TABLE {V(VCC,VEE)} =
*+({VCC1},{TPDELAY1/TPDELAY4})
*+({VCC2},{TPDELAY2/TPDELAY4})
*+({VCC3},{TPDELAY3/TPDELAY4})
*+({VCC4},{TPDELAY4/TPDELAY4})
ETPDNORM NTPDNORM VEE TABLE {V(VCC,VEE)} =
+(2,23.5)
+(4.5,11)
+(6,9)
*R1 IN N1 {RS}
G1 IN N1 VALUE = {V(IN,N1)/(V(NTPDNORM,VEE)*RS)}
RZ IN N1 10G
C1 N1 VEE {CS}
E1 N2 VEE VALUE = {0.5*(1 + SGN(V(N1,VEE) - 0.5))}
EOUT OUT VEE N2 VEE 1
.ENDS
*$
.SUBCKT LOGIC_PP_OUTPUT_HC_1i_AND_Tristate_ST IN OUT VCC VEE
* ROH1 = {(VCC1 - VOH1)/IOH1}
* ROH2 = {(VCC2 - VOH2)/IOH2}
* ROH3 = {(VCC3 - VOH3)/IOH3}
* ROH4 = {(VCC4 - VOH4)/IOH4}
* ROH5 = {(VCC5 - VOH5)/IOH5}
* ROL1 = {(VOL1)/IOL1}
* ROL2 = {(VOL2)/IOL2}
* ROL3 = {(VOL3)/IOL3}
* ROL4 = {(VOL4)/IOL4}
* ROL5 = {(VOL5)/IOL5}
*EROH NROH VEE TABLE {V(VCC,VEE)} =
*+({VCC1},{ROH1})
*+({VCC2},{ROH2})
*+({VCC3},{ROH3})
*+({VCC4},{ROH4})
*+({VCC5},{ROH5})
*EROL NROL VEE TABLE {V(VCC,VEE)} =
*+({VCC1},{ROL1})
*+({VCC2},{ROL2})
*+({VCC3},{ROL3})
*+({VCC4},{ROL4})
*+({VCC5},{ROL5})
EROH NROH VEE TABLE {V(VCC,VEE)} =
+(2,1500)
+(4.5,20)
+(6,15.3846153846154)
EROL NROL VEE TABLE {V(VCC,VEE)} =
+(2,60)
+(4.5,18)
+(6,16.9230769230769)
E1 N1 VEE VALUE = {V(VCC,VEE)*V(IN,VEE)}
GOUT N1 OUT VALUE = {V(N1,OUT)*(V(IN,VEE)/V(NROH,VEE) + (1 - V(IN,VEE))/V(NROL,VEE))}
.ENDS
*$
.SUBCKT LOGIC_OD_OUTPUT_HC_1i_AND_Tristate_ST IN OUT VCC VEE
.PARAM VCC1 = 1.65
.PARAM VCC2 = 2.3
.PARAM VCC3 = 3
.PARAM VCC4 = 3
.PARAM VCC5 = 4.5
.PARAM VOL1 = 0.45
.PARAM VOL2 = 0.3
.PARAM VOL3 = 0.4
.PARAM VOL4 = 0.55
.PARAM VOL5 = 0.55
.PARAM IOL1 = 0.004
.PARAM IOL2 = 0.008
.PARAM IOL3 = 0.016
.PARAM IOL4 = 0.024
.PARAM IOL5 = 0.032
.PARAM ROL1 = {(VOL1)/IOL1}
.PARAM ROL2 = {(VOL2)/IOL2}
.PARAM ROL3 = {(VOL3)/IOL3}
.PARAM ROL4 = {(VOL4)/IOL4}
.PARAM ROL5 = {(VOL5)/IOL5}
*EROL NROLx VEE TABLE {V(VCC,VEE)} =
*+({VCC1},{ROL1})
*+({VCC2},{ROL2})
*+({VCC4},{ROL4})
*+({VCC5},{ROL5})
EROL NROLx VEE TABLE {V(VCC,VEE)} =
+(1.65,112.5)
+(2.3,37.5)
+(3,25)
+(3,22.9166666666667)
+(4.5,17.1875)
GOUT OUT VEE VALUE = {V(OUT,VEE)*((1 - V(IN,VEE))/V(NROLx,VEE) + (1e-7)*(V(IN,VEE)))}
.ENDS
*$
.SUBCKT LOGIC_TRI_STATE_OUTPUT_HC_1i_AND_Tristate_ST IN OUT OEZ VCC VEE
.PARAM VCC1 = 4.5
.PARAM VCC2 = 5.5
.PARAM VOH1 = 4.4
.PARAM VOH2 = 3.98
.PARAM VOL1 = 0.1
.PARAM VOL2 = 0.26
.PARAM IOH1 = 0.00002
.PARAM IOH2 = 0.006
.PARAM IOL1 = 0.00002
.PARAM IOL2 = 0.006
.PARAM ROH1 = {(VCC1 - VOH1)/IOH1}
.PARAM ROH2 = {(VCC2 - VOH2)/IOH2}
.PARAM ROH3 = {(VCC3 - VOH3)/IOH3}
.PARAM ROH4 = {(VCC4 - VOH4)/IOH4}
.PARAM ROH5 = {(VCC5 - VOH5)/IOH5}
.PARAM ROL1 = {(VOL1)/IOL1}
.PARAM ROL2 = {(VOL2)/IOL2}
.PARAM ROL3 = {(VOL3)/IOL3}
.PARAM ROL4 = {(VOL4)/IOL4}
.PARAM ROL5 = {(VOL5)/IOL5}
*EROH NROH VEE TABLE {V(VCC,VEE)} =
*+({VCC1},{ROH1})
*+({VCC2},{ROH2})
*+({VCC3},{ROH3})
*+({VCC4},{ROH4})
*+({VCC5},{ROH5})
*EROL NROL VEE TABLE {V(VCC,VEE)} =
*+({VCC1},{ROL1})
*+({VCC2},{ROL2})
*+({VCC3},{ROL3})
*+({VCC4},{ROL4})
*+({VCC5},{ROL5})
EROH NROH VEE TABLE {V(VCC,VEE)} =
+(4.5,4999.99999999998)
+(5.5,253.333333333333)
EROL NROL VEE TABLE {V(VCC,VEE)} =
+(4.5,5000)
+(5.5,43.3333333333333)
EOEZ N2 VEE VALUE = {1 - V(OEZ,VEE)}
E1 N1 VEE VALUE = {V(VCC,VEE)*V(IN,VEE)*V(N2,VEE)}
GOUT N1 OUT VALUE = {V(N1,OUT)*V(N2,VEE)*(V(IN,VEE)/V(NROH,VEE) + (1 - V(IN,VEE))/V(NROL,VEE))}
LOUT N1 OUT .1n
ROUT OUT VEE 1E8
.ENDS
*$
.SUBCKT LOGIC_ICC_HC_1i_AND_Tristate_ST VCC VEE VIOUT
.PARAM ICC = 2.5e-08
.PARAM VCC_MAX = 6
.PARAM VCC_MIN = 2
*GICC VCC VEE VALUE = {ICC*V(VCC,VEE)/VCC_MAX}
GICC VCC VEE VALUE = {ICC*0.5*(1 + SGN(V(VCC,VEE) - VCC_MIN))}
*
* Floating ground at mid-rail
EGNDF GNDF 0 VALUE = {0.5*(V(VCC) + V(VEE))}
*
GOUTP VCC GNDF VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
GOUTN GNDF VEE VALUE = {V(VIOUT,VEE)*0.5*(SGN(V(VIOUT,VEE)) + ABS(SGN(V(VIOUT,VEE))))}
*
*GOUTP VCC GNDF VALUE = {IF(V(VIMON,GNDF) > 0, V(VIMON,GNDF),0)}
*GOUTN GNDF VEE VALUE = {IF(V(VIMON,GNDF) <= 0, V(VIMON,GNDF),0)}
.ENDS
*$
